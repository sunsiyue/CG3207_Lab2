----------------------------------------------------------------------------------
-- Company: NUS
-- Engineer: Rajesh Panicker
-- 
-- Create Date:   10:39:18 13/09/2014
-- Design Name: 	TOP (ALU_Test)
-- Target Devices: Nexys 4 (Artix 7 100T)
-- Tool versions: ISE 14.7
-- Description: ALU Test Wrapper
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
-- Uses uart.vhd by (c) Peter A Bennett
----------------------------------------------------------------------------------

-- NOTE : 
-- BTNC(E16) will reset both the wrapper and the ALU (Recommended)
-- BTND(V10) resets the ALU alone

-- DO NOT EDIT THIS FILE UNLESS YOU HAVE A GOOD REASON

----------------------------------------------------------------------------
-- UART Wrapper / Top Level Module
----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity TOP is
	port 
    (
	CLOCK     	: in     std_logic;
	RESET     	: in     std_logic; 
	RESET_ALU 	: in     std_logic;
	RX        	: in     std_logic;
	TX        	: out    std_logic;
	LEDS			: out 	std_logic_vector(3 downto 0); -- debug, byte counter, see UCF file for mappings
	STATE_LED	: out 	std_logic_vector(1 downto 0) -- debug, state indicator, see UCF file for mappings
    );
end TOP;

architecture RTL of TOP is
----------------------------------------------------------------------------
-- UART constants
----------------------------------------------------------------------------

constant BAUD_RATE				: positive 	:= 115200;
constant CLOCK_FREQUENCY		: positive 	:= 100000000;
constant WIDTH						: integer 	:= 32;
----------------------------------------------------------------------------
-- UART component
----------------------------------------------------------------------------
component UART is
    generic (
            BAUD_RATE           : positive;
            CLOCK_FREQUENCY     : positive
        );
    port (  -- General
            CLOCK               : in      std_logic;
            RESET               : in      std_logic;    
            DATA_STREAM_IN      : in      std_logic_vector(7 downto 0);
            DATA_STREAM_IN_STB  : in      std_logic;
            DATA_STREAM_IN_ACK  : out     std_logic;
            DATA_STREAM_OUT     : out     std_logic_vector(7 downto 0);
            DATA_STREAM_OUT_STB : out     std_logic;
            DATA_STREAM_OUT_ACK : in      std_logic;
            TX                  : out     std_logic;
            RX                  : in      std_logic
         );
end component UART;
 

----------------------------------------------------------------------------
-- UART signals
----------------------------------------------------------------------------

signal uart_data_in             : std_logic_vector(7 downto 0);
signal uart_data_out            : std_logic_vector(7 downto 0);
signal uart_data_in_stb         : std_logic;
signal uart_data_in_ack         : std_logic;
signal uart_data_out_stb        : std_logic;
signal uart_data_out_ack        : std_logic;	 

----------------------------------------------------------------------------
-- ALU component
----------------------------------------------------------------------------

component alu is
generic (width 	: integer);
Port (Clk			: in	STD_LOGIC;
		Control		: in	STD_LOGIC_VECTOR (5 downto 0);
		Operand1		: in	STD_LOGIC_VECTOR (width-1 downto 0);
		Operand2		: in	STD_LOGIC_VECTOR (width-1 downto 0);
		Result1		: out	STD_LOGIC_VECTOR (width-1 downto 0);
		Result2		: out	STD_LOGIC_VECTOR (width-1 downto 0);
		Status		: out	STD_LOGIC_VECTOR (2 downto 0); -- busy (multicycle only), overflow (add and sub), zero (sub)
		Debug			: out	STD_LOGIC_VECTOR (width-1 downto 0));		
end component alu;

----------------------------------------------------------------------------
-- ALU signals
----------------------------------------------------------------------------
 
signal	Control		: STD_LOGIC_VECTOR (5 downto 0) 			:= (others=>'0');
signal	Operand1		: STD_LOGIC_VECTOR (width-1 downto 0) 	:= (others=>'0');
signal	Operand2		: STD_LOGIC_VECTOR (width-1 downto 0) 	:= (others=>'0');
signal	Result1		: STD_LOGIC_VECTOR (width-1 downto 0) 	:= (others=>'0');
signal	Result2		: STD_LOGIC_VECTOR (width-1 downto 0) 	:= (others=>'0');
signal	Status		: STD_LOGIC_VECTOR (2 downto 0) 			:= (others=>'0');
signal	Debug			: STD_LOGIC_VECTOR (width-1 downto 0) 	:= (others=>'0');

type states is (WAITING, SENDING, PROCESSING, RECEIVING);
signal state : states := WAITING;

signal bytecounter 	: STD_LOGIC_VECTOR (4 downto 0) := (others=>'0'); -- to keep track of the bytes sent
signal cyclecounter 	: STD_LOGIC_VECTOR (15 downto 0) := (others=>'0'); -- to keep track of the cycles taken for an operation
signal storage 		: STD_LOGIC_VECTOR (114 downto 0) := (others=>'0'); --
signal uart_data_out_stb_prev : STD_LOGIC := '0';

begin

----------------------------------------------------------------------------
-- UART instantiation
----------------------------------------------------------------------------

UART1 : UART
generic map (
        BAUD_RATE           => BAUD_RATE,
        CLOCK_FREQUENCY     => CLOCK_FREQUENCY
)
port map    (  
        CLOCK               => CLOCK,
        RESET               => RESET,
        DATA_STREAM_IN      => uart_data_in,
        DATA_STREAM_IN_STB  => uart_data_in_stb,
        DATA_STREAM_IN_ACK  => uart_data_in_ack,
        DATA_STREAM_OUT     => uart_data_out,
        DATA_STREAM_OUT_STB => uart_data_out_stb,
        DATA_STREAM_OUT_ACK => uart_data_out_ack,
        TX                  => TX,
        RX                  => RX
);
 
----------------------------------------------------------------------------
-- ALU instantiation
----------------------------------------------------------------------------
 ALU1 : ALU
 generic map (width =>  width)
 port map (
		Clk => CLOCK,
		Control => Control,	
		Operand1 => Operand1,
		Operand2 => Operand2,
		Result1 => Result1,	
		Result2 => Result2,
		Status => Status,
		Debug	 => Debug
	);

Control(5) <= RESET_ALU or RESET;
LEDS <= bytecounter(3 downto 0);  --debug

UART_TOP : process (CLOCK)
begin
    if rising_edge(CLOCK) then
        if RESET = '1' then
            uart_data_in_stb        <= '0';
            uart_data_out_ack       <= '0';
            uart_data_in            <= (others => '0');
				 state 						<= WAITING;
				 Operand1 <= (others=>'0');
				 Operand2 <= (others=>'0');
				 Control(4 downto 0) <= (others=>'0');
				 uart_data_out_stb_prev <= '0';
        else
				uart_data_out_ack       <= '0';
				case state is 
					when WAITING =>
						uart_data_out_ack    <= '0';
						bytecounter <= (others=>'0');
						 if uart_data_out_stb = '1' then
							  uart_data_out_ack   <= '1';
								if uart_data_out = x"3C" then  -- '<' to begin setting
									state <= RECEIVING;	
									storage (114 downto 0) <= (others=>'0');
								end if;
						 end if;
							
					when RECEIVING =>
						uart_data_out_ack    <= '0';
						if uart_data_out_stb = '1' and uart_data_out_stb_prev = '0' then
							  uart_data_out_ack   <= '1';
							  bytecounter <= bytecounter+1;
							  case bytecounter is 
									when "00000" => storage (71 downto 64) <= uart_data_out;
									when "00001" => storage (63 downto 56) <= uart_data_out;
									when "00010" => storage (55 downto 48) <= uart_data_out;
									when "00011" => storage (47 downto 40) <= uart_data_out;
									when "00100" => storage (39 downto 32) <= uart_data_out;
									when "00101" => storage (31 downto 24) <= uart_data_out;
									when "00110" => storage (23 downto 16) <= uart_data_out;
									when "00111" => storage (15 downto 8) <= uart_data_out;
									when "01000" => storage (7 downto 0) <= uart_data_out;
									when others => 
										if uart_data_out = x"0D" then  -- '\r' to end setting, allows time to copy the buffer to inputs
											Control(4 downto 0) <= storage (68 downto 64);
											Operand1 <= storage (63 downto 32);
											Operand2 <= storage (31 downto 0);											
											state <= PROCESSING;
											cyclecounter <= x"0000";
										else -- if '\r' is not presented as expected, abort the data
											state <= WAITING;
										end if;
								end case;
						end if;
					when PROCESSING =>
						if Status(2) = '0' or cyclecounter = x"FFFF" then
							state <= SENDING;
							bytecounter <= (others=>'0');
							if Status(2) = '0' then
								storage (114 downto 112) <= '0'&Status(1 downto 0);
								storage (111 downto 96) <= cyclecounter;
								storage (95 downto 64) <= Debug;
								storage (63 downto 32) <= Result2;
								storage (31 downto 0) <= Result1;
							else   --timeout
								storage (114 downto 0) <= (114=>'1', others => '0');
							end if;
							--reset inputs immediately
							Operand1 <= (others=>'0');
							Operand2 <= (others=>'0');
							Control(4 downto 0) <= (others=>'0');
							
							uart_data_in <= x"3E";  -- > as begining of result, allows uart_data_in_ack to be checked every cycle
							uart_data_in_stb    <= '1';
						else
							cyclecounter <= cyclecounter+1;
						end if;
					
					when SENDING =>
						uart_data_in_stb <= '1';
						if uart_data_in_ack = '1' then											
							bytecounter <= bytecounter+1;
							case bytecounter is 
									 when "00000" =>uart_data_in <= "00000"& storage (114 downto 112);
									 when "00001" =>uart_data_in <= storage (111 downto 104);
									 when "00010" =>uart_data_in <= storage (103 downto 96);
									 when "00011" =>uart_data_in <= storage (95 downto 88);
									 when "00100" =>uart_data_in <= storage (87 downto 80); 
									 when "00101" =>uart_data_in <= storage (79 downto 72); 
									 when "00110" =>uart_data_in <= storage (71 downto 64); 
									 when "00111" =>uart_data_in <= storage (63 downto 56); 
									 when "01000" =>uart_data_in <= storage (55 downto 48); 
									 when "01001" =>uart_data_in <= storage (47 downto 40); 
									 when "01010" =>uart_data_in <= storage (39 downto 32); 
									 when "01011" =>uart_data_in <= storage (31 downto 24); 
									 when "01100" =>uart_data_in <= storage (23 downto 16); 
									 when "01101" =>uart_data_in <= storage (15 downto 8);
									 when "01110" =>uart_data_in <= storage (7 downto 0);
									 when "01111" =>uart_data_in <= x"0D"; --'\r' as end of result
									 when others => 
												state <= WAITING;
												uart_data_in_stb    <= '0';
							end case;
						end if;
				end case; 
        end if;
			uart_data_out_stb_prev <= uart_data_out_stb;
    end if;
end process;
 
state_indicator : process(state)
begin
	case state is
		when WAITING 		=> 	STATE_LED <= "00";
		when RECEIVING 	=> 	STATE_LED <= "01";
		when PROCESSING 	=> 	STATE_LED <= "10";
		when SENDING 		=> 	STATE_LED <= "11";  
	end case;
end process;

end RTL;

